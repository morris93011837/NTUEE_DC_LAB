
module rsa_qsys (
	clk_clk,
	reset_reset_n,
	altpll_100k_clk,
	altpll_12m_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		altpll_100k_clk;
	output		altpll_12m_clk;
endmodule
